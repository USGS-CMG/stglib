version https://git-lfs.github.com/spec/v1
oid sha256:0c58180ae2d90370bfd9de6178c258fd0bba33319787b9581c087a5751521f6e
size 869850

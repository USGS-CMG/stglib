version https://git-lfs.github.com/spec/v1
oid sha256:016f4c2cff24a54e8d5e573edadea6b8610ebc38df587e37c7f60326d376791d
size 150
